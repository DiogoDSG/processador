library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ram_tb is
end entity;

architecture a_ram_tb of ram_tb is
    component ram
        port(  
            clk : in std_logic;
            address : in unsigned(6 downto 0);
            wr_en : in std_logic;
            data_in : in unsigned(15 downto 0);
            data_out : out unsigned(15 downto 0)
        ); 
    end component;

    constant period_time: time := 100 ns;
    signal wr_en, clk: std_logic;
    signal data_in, data_out: unsigned(15 downto 0);
    signal finished: std_logic := '0';
    signal address: unsigned(6 downto 0);
    begin
        uut: ram port map(
            clk => clk,
            address => address,
            wr_en => wr_en,
            data_in => data_in,
            data_out => data_out
        );

    sim_time_proc: process
    begin
        wait for 100 us;
        finished <= '1';
        wait;
    end process;

    clk_global: process
    begin
        while finished /= '1' loop
            clk <= '1';
            wait for period_time / 2;
            clk <= '0';
            wait for period_time / 2;
        end loop;
        wait;
    end process;


    process
    begin
        wr_en <= '1';
        wait for period_time;
        data_in <= "0000000000000000";
        address <= "0000000";
        wait for period_time;
        data_in <= "0000000000000001";
        address <= "0000001";
        wait for period_time;
        data_in <= "0000000000000010";
        address <= "0000010";
        wait for period_time;
        data_in <= "0000000000000011";
        address <= "0000011";
        wait for period_time;
        data_in <= "0000000000000100";
        address <= "0000100";
        wait for period_time;
        data_in <= "0000000000000101";
        address <= "0000101";
        wait for period_time;
        data_in <= "0000000000000110";
        address <= "0000110";
        wait for period_time;
        data_in <= "0000000000000111";
        address <= "0000111";
        wait for period_time;
        data_in <= "0000000000001000";
        address <= "0001000";
        wait for period_time;
        data_in <= "0000000000001001";
        address <= "0001001";
        wait for period_time;
        data_in <= "0000000000001010";
        address <= "0001010";
        wait for period_time;
        data_in <= "0000000000001011";
        address <= "0001011";
        wait for period_time;
        data_in <= "0000000000001100";
        address <= "0001100";
        wait for period_time;
        data_in <= "0000000000001101";
        address <= "0001101";
        wait for period_time;
        data_in <= "0000000000001110";
        address <= "0001110";
        wait for period_time;
        data_in <= "0000000000001111";
        address <= "0001111";
        wait for period_time;
        data_in <= "0000000000010000";
        address <= "0010000";
        wait for period_time;
        data_in <= "0000000000010001";
        address <= "0010001";
        wait for period_time;
        data_in <= "0000000000010010";
        address <= "0010010";
        wait for period_time;
        data_in <= "0000000000010011";
        address <= "0010011";
        wait for period_time;
        data_in <= "0000000000010100";
        address <= "0010100";
        wait for period_time;
        data_in <= "0000000000010101";
        address <= "0010101";
        wait for period_time;
        data_in <= "0000000000010110";
        address <= "0010110";
        wait for period_time;
        data_in <= "0000000000010111";
        address <= "0010111";
        wait for period_time;
        data_in <= "0000000000011000";
        address <= "0011000";
        wait for period_time;
        data_in <= "0000000000011001";
        address <= "0011001";
        wait for period_time;
        data_in <= "0000000000011010";
        address <= "0011010";
        wait for period_time;
        data_in <= "0000000000011011";
        address <= "0011011";
        wait for period_time;
        data_in <= "0000000000011100";
        address <= "0011100";
        wait for period_time;
        data_in <= "0000000000011101";
        address <= "0011101";
        wait for period_time;
        data_in <= "0000000000011110";
        address <= "0011110";
        wait for period_time;
        data_in <= "0000000000011111";
        address <= "0011111";
        wait for period_time;
        data_in <= "0000000000100000";
        address <= "0100000";
        wait for period_time;
        data_in <= "0000000000100001";
        address <= "0100001";
        wait for period_time;
        data_in <= "0000000000100010";
        address <= "0100010";
        wait for period_time;
        data_in <= "0000000000100011";
        address <= "0100011";
        wait for period_time;
        data_in <= "0000000000100100";
        address <= "0100100";
        wait for period_time;
        data_in <= "0000000000100101";
        address <= "0100101";
        wait for period_time;
        data_in <= "0000000000100110";
        address <= "0100110";
        wait for period_time;
        data_in <= "0000000000100111";
        address <= "0100111";
        wait for period_time;
        data_in <= "0000000000101000";
        address <= "0101000";
        wait for period_time;
        data_in <= "0000000000101001";
        address <= "0101001";
        wait for period_time;
        data_in <= "0000000000101010";
        address <= "0101010";
        wait for period_time;
        data_in <= "0000000000101011";
        address <= "0101011";
        wait for period_time;
        data_in <= "0000000000101100";
        address <= "0101100";
        wait for period_time;
        data_in <= "0000000000101101";
        address <= "0101101";
        wait for period_time;
        data_in <= "0000000000101110";
        address <= "0101110";
        wait for period_time;
        data_in <= "0000000000101111";
        address <= "0101111";
        wait for period_time;
        data_in <= "0000000000110000";
        address <= "0110000";
        wait for period_time;
        data_in <= "0000000000110001";
        address <= "0110001";
        wait for period_time;
        data_in <= "0000000000110010";
        address <= "0110010";
        wait for period_time;
        data_in <= "0000000000110011";
        address <= "0110011";
        wait for period_time;
        data_in <= "0000000000110100";
        address <= "0110100";
        wait for period_time;
        data_in <= "0000000000110101";
        address <= "0110101";
        wait for period_time;
        data_in <= "0000000000110110";
        address <= "0110110";
        wait for period_time;
        data_in <= "0000000000110111";
        address <= "0110111";
        wait for period_time;
        data_in <= "0000000000111000";
        address <= "0111000";
        wait for period_time;
        data_in <= "0000000000111001";
        address <= "0111001";
        wait for period_time;
        data_in <= "0000000000111010";
        address <= "0111010";
        wait for period_time;
        data_in <= "0000000000111011";
        address <= "0111011";
        wait for period_time;
        data_in <= "0000000000111100";
        address <= "0111100";
        wait for period_time;
        data_in <= "0000000000111101";
        address <= "0111101";
        wait for period_time;
        data_in <= "0000000000111110";
        address <= "0111110";
        wait for period_time;
        data_in <= "0000000000111111";
        address <= "0111111";
        wait for period_time;
        data_in <= "0000000001000000";
        address <= "1000000";
        wait for period_time;
        data_in <= "0000000001000001";
        address <= "1000001";
        wait for period_time;
        data_in <= "0000000001000010";
        address <= "1000010";
        wait for period_time;
        data_in <= "0000000001000011";
        address <= "1000011";
        wait for period_time;
        data_in <= "0000000001000100";
        address <= "1000100";
        wait for period_time;
        data_in <= "0000000001000101";
        address <= "1000101";
        wait for period_time;
        data_in <= "0000000001000110";
        address <= "1000110";
        wait for period_time;
        data_in <= "0000000001000111";
        address <= "1000111";
        wait for period_time;
        data_in <= "0000000001001000";
        address <= "1001000";
        wait for period_time;
        data_in <= "0000000001001001";
        address <= "1001001";
        wait for period_time;
        data_in <= "0000000001001010";
        address <= "1001010";
        wait for period_time;
        data_in <= "0000000001001011";
        address <= "1001011";
        wait for period_time;
        data_in <= "0000000001001100";
        address <= "1001100";
        wait for period_time;
        data_in <= "0000000001001101";
        address <= "1001101";
        wait for period_time;
        data_in <= "0000000001001110";
        address <= "1001110";
        wait for period_time;
        data_in <= "0000000001001111";
        address <= "1001111";
        wait for period_time;
        data_in <= "0000000001010000";
        address <= "1010000";
        wait for period_time;
        data_in <= "0000000001010001";
        address <= "1010001";
        wait for period_time;
        data_in <= "0000000001010010";
        address <= "1010010";
        wait for period_time;
        data_in <= "0000000001010011";
        address <= "1010011";
        wait for period_time;
        data_in <= "0000000001010100";
        address <= "1010100";
        wait for period_time;
        data_in <= "0000000001010101";
        address <= "1010101";
        wait for period_time;
        data_in <= "0000000001010110";
        address <= "1010110";
        wait for period_time;
        data_in <= "0000000001010111";
        address <= "1010111";
        wait for period_time;
        data_in <= "0000000001011000";
        address <= "1011000";
        wait for period_time;
        data_in <= "0000000001011001";
        address <= "1011001";
        wait for period_time;
        data_in <= "0000000001011010";
        address <= "1011010";
        wait for period_time;
        data_in <= "0000000001011011";
        address <= "1011011";
        wait for period_time;
        data_in <= "0000000001011100";
        address <= "1011100";
        wait for period_time;
        data_in <= "0000000001011101";
        address <= "1011101";
        wait for period_time;
        data_in <= "0000000001011110";
        address <= "1011110";
        wait for period_time;
        data_in <= "0000000001011111";
        address <= "1011111";
        wait for period_time;
        data_in <= "0000000001100000";
        address <= "1100000";
        wait for period_time;
        data_in <= "0000000001100001";
        address <= "1100001";
        wait for period_time;
        data_in <= "0000000001100010";
        address <= "1100010";
        wait for period_time;
        data_in <= "0000000001100011";
        address <= "1100011";
        wait for period_time;
        data_in <= "0000000001100100";
        address <= "1100100";
        wait for period_time;
        data_in <= "0000000001100101";
        address <= "1100101";
        wait for period_time;
        data_in <= "0000000001100110";
        address <= "1100110";
        wait for period_time;
        data_in <= "0000000001100111";
        address <= "1100111";
        wait for period_time;
        data_in <= "0000000001101000";
        address <= "1101000";
        wait for period_time;
        data_in <= "0000000001101001";
        address <= "1101001";
        wait for period_time;
        data_in <= "0000000001101010";
        address <= "1101010";
        wait for period_time;
        data_in <= "0000000001101011";
        address <= "1101011";
        wait for period_time;
        data_in <= "0000000001101100";
        address <= "1101100";
        wait for period_time;
        data_in <= "0000000001101101";
        address <= "1101101";
        wait for period_time;
        data_in <= "0000000001101110";
        address <= "1101110";
        wait for period_time;
        data_in <= "0000000001101111";
        address <= "1101111";
        wait for period_time;
        data_in <= "0000000001110000";
        address <= "1110000";
        wait for period_time;
        data_in <= "0000000001110001";
        address <= "1110001";
        wait for period_time;
        data_in <= "0000000001110010";
        address <= "1110010";
        wait for period_time;
        data_in <= "0000000001110011";
        address <= "1110011";
        wait for period_time;
        data_in <= "0000000001110100";
        address <= "1110100";
        wait for period_time;
        data_in <= "0000000001110101";
        address <= "1110101";
        wait for period_time;
        data_in <= "0000000001110110";
        address <= "1110110";
        wait for period_time;
        data_in <= "0000000001110111";
        address <= "1110111";
        wait for period_time;
        data_in <= "0000000001111000";
        address <= "1111000";
        wait for period_time;
        data_in <= "0000000001111001";
        address <= "1111001";
        wait for period_time;
        data_in <= "0000000001111010";
        address <= "1111010";
        wait for period_time;
        data_in <= "0000000001111011";
        address <= "1111011";
        wait for period_time;
        data_in <= "0000000001111100";
        address <= "1111100";
        wait for period_time;
        data_in <= "0000000001111101";
        address <= "1111101";
        wait for period_time;
        data_in <= "0000000001111110";
        address <= "1111110";
        wait for period_time;
        data_in <= "0000000001111111";
        address <= "1111111";
        wait for period_time;
        wr_en <= '0';
        data_in <= "0011100000000000";
        address <= "0000001";
        wait for period_time;
        address <= "0000000";
        wait for period_time;
        address <= "0000001";
        wait;
    end process;
end architecture;