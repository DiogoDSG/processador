
library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 
entity rom is   
    port(         
    address: in unsigned(6 downto 0);         
    data: out unsigned(13 downto 0)); 
end entity; 
architecture a_rom of rom is type mem is array (0 to 127) of unsigned(13 downto 0);   
constant rom_content : mem := (
    0 => "01100010000010",
    1 => "01100100000100",
    2 => "01011110010000",
    3 => "01101010000111",
    4 => "00011111110100",
    5 => "00000000000000",
    6 => "01010111110000",
    7 => "00000000000000",
    8 => "01101110000000",
    9 => "00000000000000",
    10 => "01011111010000",
    11 => "00000000000000",
    12 => "00101111110010",
    13 => "00000000000000",
    14 => "01011001110000",
    15 => "00000000000000",
    16 => "01101110000000",
    17 => "00000000000000",
    18 => "11110000000000",
    19 => "00000000000000",



    -- 0  => "01100010000010",
    -- 1  => "01100100000100",  
    -- 2  => "01101010000111",          
    -- 3  => "00010110010100",      
    -- 4  => "00101001010010",  
    -- 5  => "01011100110000",
    -- 6  => "00000000000000",
    -- 6  => "11110000000000",    
    -- 4  => "10000000000000",      
    -- 5  => "00000000001000",      
    -- 6  => "11110000000000",      
    -- 7  => "00000000001000",      
    -- 8  => "00000000001000",      
    -- 9  => "00000000000000",      
    -- 10 => "00000000000000",
    -- abaixo: casos omissos => (zero em todos os bits)      
    others => (others=>'0'));    
    begin
    data <= rom_content(to_integer(address));      
 
end architecture;