
library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 
entity rom is   
    port(         
    address: in unsigned(6 downto 0);         
    data: out unsigned(13 downto 0)); 
end entity; 
architecture a_rom of rom is type mem is array (0 to 127) of unsigned(13 downto 0);   
constant rom_content : mem := (
    0 => "01010110000001",
	1 => "01011000000001",
	2 => "01011110110000",
	3 => "00000000000000",
	4 => "00000000000000",
	5 => "00000000000000",
	6 => "00011000000000",
	7 => "00000000000000",
	8 => "00000000000000",
	9 => "00000000000000",
	10 => "01011001110000",
	11 => "00000000000000",
	12 => "00000000000000",
	13 => "00000000000000",
	14 => "01011110110000",
	15 => "01010010000011",
	16 => "00000000000000",
	17 => "00000000000000",
	18 => "00000000000000",
	19 => "00010010000000",
	20 => "00000000000000",
	21 => "00000000000000",
	22 => "00000000000000",
	23 => "01010111110000",
	24 => "01011100111101",
	25 => "01011110110000",
	26 => "00000000000000",
	27 => "00000000000000",
	28 => "00000000000000",
	29 => "00101100000000",
	30 => "11100000000010",
	
    others => (others=>'0'));    
    begin
    data <= rom_content(to_integer(address));      
 
end architecture;
