
library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 
entity rom is   
    port(         
    address: in unsigned(6 downto 0);         
    data: out unsigned(13 downto 0)); 
end entity; 
architecture a_rom of rom is type mem is array (0 to 127) of unsigned(13 downto 0);   
constant rom_content : mem := (
    0 => "01011110000011",
	1 => "01010010000011",
	2 => "01110001110000",
	3 => "00010000000011",
	4 => "00110001000011",
	5 => "11100000000010",
	6 => "01011110010000",
	7 => "00010000000011",
	8 => "00110000000000",
	9 => "11000000000110",
	10 => "01010011110000",
	11 => "00010010000000",
	12 => "01010101110000",
	13 => "01011110000001",
	14 => "01110000100000",
	15 => "01011110100000",
	16 => "00110001000011",
	17 => "11100000001011",
	18 => "01011110010000",
	19 => "00110001000011",
	20 => "11100000000110",
	21 => "01010110000011",
	22 => "01100000110000",
	23 => "01011001110000",
	24 => "01011110110000",
	25 => "00010000000011",
	26 => "01010111110000",
	27 => "00110001000011",
	28 => "11100000010110",
	
    others => (others=>'0'));    
    begin
    data <= rom_content(to_integer(address));      
 
end architecture;
